-- Vhdl test bench created from schematic C:\Users\160544C\Documents\WorkSpace\Lab_4\Decoder_3_8.sch - Thu Sep 14 13:54:21 2017
--
-- Notes: 
-- 1) This testbench template has been automatically generated using types
-- std_logic and std_logic_vector for the ports of the unit under test.
-- Xilinx recommends that these types always be used for the top-level
-- I/O of a design in order to guarantee that the testbench will bind
-- correctly to the timing (post-route) simulation model.
-- 2) To use this template as your testbench, change the filename to any
-- name of your choice with the extension .vhd, and use the "Source->Add"
-- menu in Project Navigator to import the testbench. Then
-- edit the user defined section below, adding code to generate the 
-- stimulus for your design.
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
LIBRARY UNISIM;
USE UNISIM.Vcomponents.ALL;
ENTITY Decoder_3_8_Decoder_3_8_sch_tb IS
END Decoder_3_8_Decoder_3_8_sch_tb;
ARCHITECTURE behavioral OF Decoder_3_8_Decoder_3_8_sch_tb IS 

   COMPONENT Decoder_3_8
   PORT( );
   END COMPONENT;


BEGIN

   UUT: Decoder_3_8 PORT MAP(
		
   );

-- *** Test Bench - User Defined Section ***
   tb : PROCESS
   BEGIN
      WAIT; -- will wait forever
   END PROCESS;
-- *** End Test Bench - User Defined Section ***

END;
